module toplevel(input btnC, input btnU, input btnL, input btnR, input btnD, input swt, input clk, output [3:0] JC);

   main main_module(btnC, btnU, btnL, btnR, btnD, swt, clk, ,);
   //TODO, include the music decoder
   //make the output thing 

endmodule //ligma
