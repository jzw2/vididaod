module toplevel(input btnC, input btnU, input btnL, input btnR, input btnD, input swt, input clk, output y);

   main main_module(btC, btU, btnL, btnR, btnD, swt, clk, ,);
   //make the output thing 

endmodule; //ligma
